** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/CMOS_Char/Ron_test.sch
**.subckt Ron_test
XM1 Vd Vg GND GND sg13_hv_nmos w={W} l=0.45u ng=1 m=1
Vg Vg GND 3.3
Vd Vd GND 3.3
**** begin user architecture code



.control
save all
+ @n.xm1.nsg13_hv_nmos[gds]
op
let rds =1/@n.xm1.nsg13_hv_nmos[gds]
print rds
.endc



.lib cornerMOShv.lib mos_tt




.param W = 1.0u
.param Vdd = 3.3


**** end user architecture code
**.ends
.GLOBAL GND
.end
