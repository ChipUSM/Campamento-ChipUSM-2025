** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/TRAN_NOT.sch
**.subckt TRAN_NOT VOUT VIN
*.iopin VOUT
*.iopin VIN
x1 VDD VIN VOUT GND NOT
C1 VOUT GND 25f m=1
V1 VDD GND 3.3
**** begin user architecture code


.lib cornerMOShv.lib mos_tt
.lib cornerMOSlv.lib mos_tt
*.lib cornerMOShv.lib mos_ff
*.lib cornerMOSlv.lib mos_ff
*.lib cornerMOShv.lib mos_ss
*.lib cornerMOSlv.lib mos_ss
*.lib cornerMOShv.lib mos_sf
*.lib cornerMOSlv.lib mos_sf
*.lib cornerMOShv.lib mos_fs
*.lib cornerMOSlv.lib mos_fs

*.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/diodes.lib



vin VIN 0 PULSE(0 3.3 1ns 0ns 0ns 2ns 4ns)

.control
save all
***********************************************
* SIMULACION DE 10 NANO DE DURACION, CON MEDICIONES CADA 100 PICO
tran 100ps 10ns

**********************************************

plot V(VIN) v(VOUT)

**********************************************
*COMANDOS PARA MEDIR EL TIEMPO DE PROPAGACIÓN DE LA COMPUERTA

meas tran tpLH_in FIND time WHEN v(VIN)=1.65 TD=0 FALL=1
meas tran tpLH_fin FIND time WHEN v(VOUT)=1.65 TD=0 RISE=1
meas tran tpHL_in FIND time WHEN v(VIN)=1.65 TD=0 RISE=1
meas tran tpHL_fin FIND time WHEN v(VOUT)=1.65 TD=0 FALL=1
print tpHL_fin - tpHL_in
print tpLH_fin - tpLH_in
**********************************************
.endc


**** end user architecture code
**.ends

* expanding   symbol:  ../LogicGates/NOT.sym # of pins=4
** sym_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/NOT.sym
** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/NOT.sch
.subckt NOT VDD Vin Vout GND
*.ipin VDD
*.ipin Vin
*.ipin GND
*.opin Vout
XM3 GND Vin Vout GND sg13_hv_nmos w=1.0u l=0.45u ng=1 m=1
XM4 Vout Vin VDD VDD sg13_hv_pmos w=2.72u l=0.45u ng=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
