** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/TB_NAND.sch
**.subckt TB_NAND
V1 Vdd GND {Vdd}
C1 out GND 1f m=1
x1 Vdd A B out GND NAND
V2 A GND PULSE(0 {Vdd} {T/2} {T/200} {T/200} {T/2} {T})
V3 B GND PULSE(0 {Vdd} {T} {T/200} {T/200} {T} {2*T})
**** begin user architecture code



.control
save all

tran 10p 10n

meas tran Propagacion_Low_High TRIG v(a) VAL=0.6 RISE=2 TARG v(out) VAL=0.6 FALL=1
plot v(A) v(B) (v(out) + 1.2)
.endc





.lib cornerMOSlv.lib mos_tt



.param T = 2n
.param Vdd = 1.2
.param W_n = 1u
.param W_p = 1u


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/NAND.sym # of pins=5
** sym_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/NAND.sym
** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/LogicGates/NAND.sch
.subckt NAND Vdd A B F Vss
*.ipin Vss
*.ipin A
*.ipin B
*.ipin Vdd
*.opin F
XM1 F B net1 Vss sg13_lv_nmos w={W_n} l=0.13u ng=1 m=1
XM2 net1 A Vss Vss sg13_lv_nmos w={W_n} l=0.13u ng=1 m=1
XM3 F B Vdd Vdd sg13_lv_pmos w={W_p} l=0.13u ng=1 m=1
XM4 F A Vdd Vdd sg13_lv_pmos w={W_n} l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
