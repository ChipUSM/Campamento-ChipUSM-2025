** sch_path: /foss/designs/Campamento-ChipUSM-2025/xschem/CMOS_Char/Vgs_HvMOS.sch
**.subckt Vgs_HvMOS
XM1 Vd Vg GND GND sg13_hv_nmos w=10u l=0.45u ng=1 m=1
Vg Vg GND 3.3
Vd Vd GND 3.3
XM2 Vd Vg GND GND sg13_hv_nmos w=10u l=0.45u ng=2 m=1
XM3 Vd Vg GND GND sg13_hv_nmos w=5u l=0.45u ng=1 m=2
**** begin user architecture code



.control

*** ALMACENAR DATOS Y CORRER SIMULACION

save all
+ @n.xm1.nsg13_hv_nmos[vgs]
+ @n.xm1.nsg13_hv_nmos[ids]
+ @n.xm1.nsg13_hv_nmos[gm]
+ @n.xm2.nsg13_hv_nmos[vgs]
+ @n.xm2.nsg13_hv_nmos[ids]
+ @n.xm2.nsg13_hv_nmos[gm]
+ @n.xm3.nsg13_hv_nmos[vgs]
+ @n.xm3.nsg13_hv_nmos[ids]
+ @n.xm3.nsg13_hv_nmos[gm]

dc Vg 0 3.3 0.01

*** GUARDAR DATOS COMO VARIABLES Y GRAFICAR

let vgs1 = @n.xm1.nsg13_hv_nmos[vgs]
let ids1 = @n.xm1.nsg13_hv_nmos[ids]
let gm1 = @n.xm1.nsg13_hv_nmos[gm]

let vgs2 = @n.xm2.nsg13_hv_nmos[vgs]
let ids2 = @n.xm2.nsg13_hv_nmos[ids]
let gm1 = @n.xm2.nsg13_hv_nmos[gm]


let vgs3 = @n.xm3.nsg13_hv_nmos[vgs]
let ids3 = @n.xm3.nsg13_hv_nmos[ids]
let gm3 = @n.xm3.nsg13_hv_nmos[gm]

plot ids1 vs vgs1
plot ids2 vs vgs2
plot ids3 vs vgs3

plot gm1 vs vgs1
print ids1[330]
print ids2[330]
print ids3[330]
.endc



.lib cornerMOShv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
